//  ###########################################################################
//
//  Licensed to the Apache Software Foundation (ASF) under one
//  or more contributor license agreements.  See the NOTICE file
//  distributed with this work for additional information
//  regarding copyright ownership.  The ASF licenses this file
//  to you under the Apache License, Version 2.0 (the
//  "License"); you may not use this file except in compliance
//  with the License.  You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing,
//  software distributed under the License is distributed on an
//  "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
//  KIND, either express or implied.  See the License for the
//  specific language governing permissions and limitations
//  under the License.
//  
//  ###########################################################################

`ifndef AXI4_TOP_SV
`define AXI4_TOP_SV

//-----------------------------------------------------------------------------
//Module : axi4_top
//Description : 
//Top module to generate the clock frequency and invoking the test cases.
//-----------------------------------------------------------------------------

module top;

bit clock;

axi_if i_f(clock);

//Clock Generation
always 
  #20 clock = ~clock;

//Invoking Test cases
initial begin
  uvm_config_db #(virtual axi_if)::set(null,"*","vif",i_f);
  run_test("base_test"); 
end

endmodule

`endif

//----E.O.F------
